`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.02.2024 22:48:33
// Design Name: 
// Module Name: alu_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu_tb();
reg [31:0]A,B;
wire [31:0]out1, out2, out3;
wire out4;
reg o;
alu_top alu1(A,B,o,out1, out2, out3, out4);



initial
begin
 A = 32'b0_10000001_00000000000000000000000;
B = 32'b0_10000000_00000000000000000000000; o = 1'b0;
#10 A = 32'b0_10000010_01000000000000000000000;
B= 32'b1_10000000_00000000000000000000000; o = 1'b0;
#10 A = 32'b0_10000001_11000000000000000000000;
B= 32'b0_10000000_00000000000000000000000; o = 1'b1;
#10 A = 32'b0_10000010_10011100110011001100110;
B= 32'b1_10000010_00100110011001100110011; o = 1'b0;
#10 A = 32'b1_10000001_01011001100110011001101; 
B= 32'b0_10000000_00100110011001100110011; o = 1'b0;
#10 $stop;

end

endmodule


